MACRO C0
     SIZE 4302 BY 2223 ;
END C0
MACRO C1
     SIZE 10418 BY 3815 ;
END C1
MACRO C2
     SIZE 8447 BY 3056 ;
END C2
MACRO C3
     SIZE 11393 BY 2149 ;
END C3
MACRO C4
     SIZE 11313 BY 6449 ;
END C4
